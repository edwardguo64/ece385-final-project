module Sprite(		
    output logic [4:0][28:0][3:0] score_letters,
	output logic [4:0][28:0][3:0] level_letters,
	output logic [4:0][22:0][3:0] line_letters,
    output logic [4:0][4:0][3:0] zero,
    output logic [4:0][4:0][3:0] one,
    output logic [4:0][4:0][3:0] two,
    output logic [4:0][4:0][3:0] three,
    output logic [4:0][4:0][3:0] four,
    output logic [4:0][4:0][3:0] five,
    output logic [4:0][4:0][3:0] six,
    output logic [4:0][4:0][3:0] seven,
    output logic [4:0][4:0][3:0] eight,
    output logic [4:0][4:0][3:0] nine,
	output logic [13:0][78:0][3:0] gameover_text,
	output logic [13:0][57:0][3:0] Game_Start,
    output logic [4:0][90:0][3:0] press_start,
    output logic [4:0][112:0][3:0] play_again,
    output logic [4:0][46:0][3:0] high_score,
    output logic [4:0][46:0][3:0] your_score
);

    always_comb
    begin
		Game_Start = '{
            '{1,1,1,1,1,1,1,1,1,0,2,2,2,2,2,2,2,2,0,3,3,3,3,3,3,3,3,3,0,4,4,4,4,4,4,4,4,0,0,0,0,0,5,5,5,0,0,0,0,1,1,1,1,1,1,1,1,1},
            '{1,1,1,1,1,1,1,1,1,0,2,2,2,2,2,2,2,2,0,3,3,3,3,3,3,3,3,3,0,4,4,4,4,4,4,4,4,0,0,0,0,0,5,5,5,0,0,0,0,1,1,1,1,1,1,1,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,0,4,4,0,0,0,0,5,5,5,0,0,0,0,1,1,0,0,0,0,0,0,0},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,0,4,4,0,0,0,0,5,5,5,0,0,0,0,1,1,0,0,0,0,0,0,0},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,0,4,4,0,0,0,0,5,5,5,0,0,0,0,1,1,0,0,0,0,0,0,0},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,0,4,4,0,0,0,0,5,5,5,0,0,0,0,1,1,0,0,0,0,0,0,0},
            '{0,0,0,1,1,1,0,0,0,0,2,2,2,2,2,2,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,4,4,4,4,4,4,0,0,0,0,0,5,5,5,0,0,0,0,1,1,1,1,1,1,1,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,2,2,2,2,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,4,4,4,4,4,4,0,0,0,0,0,5,5,5,0,0,0,0,1,1,1,1,1,1,1,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,4,4,0,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0,0,0,0,0,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,4,4,0,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0,0,0,0,0,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,4,4,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0,0,0,0,0,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,4,4,0,0,0,0,0,5,5,5,0,0,0,0,0,0,0,0,0,0,0,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,2,2,2,2,2,2,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,0,4,4,0,0,0,0,5,5,5,0,0,0,0,1,1,1,1,1,1,1,1,1},
            '{0,0,0,1,1,1,0,0,0,0,2,2,2,2,2,2,2,2,0,0,0,0,3,3,3,0,0,0,0,4,4,0,0,0,0,0,4,4,0,0,0,0,5,5,5,0,0,0,0,1,1,1,1,1,1,1,1,1}
		};
        
        press_start = '{
            '{1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,0,0,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,1,1,1,0,0,1,1,0,0,1,1,1,1,0,1,1,1,1,0},
            '{1,0,0,1,0,1,0,0,1,0,1,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,1,1,0,1,0,0,1,1,0,0,1,0,0,0,0,1,0,0,1,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,1,0,0,0,0,0,1,1,0,0,1,0,0,1,0,1,0,0,1,0,0,1,1,0,0},
            '{1,1,1,1,0,1,1,1,1,0,1,1,1,0,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,0,0,1,1,1,1,0,0,1,1,0,0,1,1,1,0,0,1,1,1,1,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,1,1,1,1,0,0,1,1,0,0,1,1,1,1,0,1,1,1,1,0,0,1,1,0,0},
            '{1,0,0,0,0,1,0,1,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,1,0,0,0,0,1,0,1,1,0,0,1,1,0,0,1,0,0,0,0,1,0,1,0,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,0,0,0,1,0,0,1,1,0,0,1,0,0,1,0,1,0,1,0,0,0,1,1,0,0},
            '{1,0,0,0,0,1,0,0,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,0,0,1,0,0,1,1,0,0,1,1,1,1,0,1,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1,0,0,0,1,1,1,1,0,0,1,1,0,0,1,0,0,1,0,1,0,0,1,0,0,1,1,0,0}
        };
		  
		gameover_text  =  '{
            '{0,1,1,1,1,1,1,0,0,0,0,0,0,2,2,2,0,0,0,0,3,3,0,0,0,0,0,3,3,0,4,4,4,4,4,4,4,4,0,0,5,5,5,5,5,5,5,0,0,1,1,0,0,0,0,0,1,1,0,2,2,2,2,2,2,2,2,0,3,3,3,3,3,3,3,3,0,0,0},
            '{0,1,1,1,1,1,1,0,0,0,0,0,0,2,2,2,0,0,0,0,3,3,0,0,0,0,0,3,3,0,4,4,4,4,4,4,4,4,0,0,5,5,5,5,5,5,5,0,0,1,1,0,0,0,0,0,1,1,0,2,2,2,2,2,2,2,2,0,3,3,3,3,3,3,3,3,0,0,0},
            '{1,1,0,0,0,0,1,1,0,0,0,0,2,2,0,2,2,0,0,0,3,3,3,0,0,0,3,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,1,1,0,0,0,0,0,1,1,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,0,0,3,3,0,0},
            '{1,1,0,0,0,0,1,1,0,0,0,0,2,2,0,2,2,0,0,0,3,3,3,0,0,0,3,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,1,1,0,0,0,0,0,1,1,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,0,0,3,3,0,0},
            '{1,1,0,0,0,0,0,0,0,0,0,2,2,0,0,0,2,2,0,0,3,3,3,3,0,3,3,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,1,1,0,0,0,0,0,1,1,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,0,0,3,3,0,0},
            '{1,1,0,0,0,0,0,0,0,0,0,2,2,0,0,0,2,2,0,0,3,3,3,3,0,3,3,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,1,1,0,0,0,0,0,1,1,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,0,0,3,3,0,0},
            '{1,1,0,0,0,1,1,1,1,0,2,2,0,0,0,0,0,2,2,0,3,3,0,3,3,3,0,3,3,0,4,4,4,4,4,4,0,0,0,5,5,0,0,0,0,0,5,5,0,1,1,0,0,0,0,0,1,1,0,2,2,2,2,2,2,0,0,0,3,3,3,3,3,3,3,3,0,0,0},
            '{1,1,0,0,0,1,1,1,1,0,2,2,0,0,0,0,0,2,2,0,3,3,0,3,3,3,0,3,3,0,4,4,4,4,4,4,0,0,0,5,5,0,0,0,0,0,5,5,0,1,1,0,0,0,0,0,1,1,0,2,2,2,2,2,2,0,0,0,3,3,3,3,3,3,3,3,0,0,0},
            '{1,1,0,0,0,0,1,1,0,0,2,2,2,2,2,2,2,2,2,0,3,3,0,0,0,0,0,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,0,1,1,0,0,0,1,1,0,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,3,3,0,0,0,0},
            '{1,1,0,0,0,0,1,1,0,0,2,2,2,2,2,2,2,2,2,0,3,3,0,0,0,0,0,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,0,1,1,0,0,0,1,1,0,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,3,3,0,0,0,0},
            '{1,1,0,0,0,0,1,1,0,0,2,2,0,0,0,0,0,2,2,0,3,3,0,0,0,0,0,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,0,0,1,1,0,1,1,0,0,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,0,3,3,0,0,0},
            '{1,1,0,0,0,0,1,1,0,0,2,2,0,0,0,0,0,2,2,0,3,3,0,0,0,0,0,3,3,0,4,4,0,0,0,0,0,0,0,5,5,0,0,0,0,0,5,5,0,0,0,1,1,0,1,1,0,0,0,2,2,0,0,0,0,0,0,0,3,3,0,0,0,0,3,3,0,0,0},
            '{0,1,1,1,1,1,1,0,0,0,2,2,0,0,0,0,0,2,2,0,3,3,0,0,0,0,0,3,3,0,4,4,4,4,4,4,4,4,0,0,5,5,5,5,5,5,5,0,0,0,0,0,1,1,1,0,0,0,0,2,2,2,2,2,2,2,2,0,3,3,0,0,0,0,0,3,3,0,0},
            '{0,1,1,1,1,1,1,0,0,0,2,2,0,0,0,0,0,2,2,0,3,3,0,0,0,0,0,3,3,0,4,4,4,4,4,4,4,4,0,0,5,5,5,5,5,5,5,0,0,0,0,0,1,1,1,0,0,0,0,2,2,2,2,2,2,2,2,0,3,3,0,0,0,0,0,3,3,0,0}
        };
        
        play_again = '{
            '{1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,0,0,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,0,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,0,0,1,0,0,1,0},
            '{1,0,0,1,0,1,0,0,1,0,1,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,1,1,0,1,0,0,1,1,0,0,1,0,0,0,0,1,0,0,1,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,1,0,0,1,0,1,0,0,0,0,1,0,0,1,0,1,0,0,1,0,0,0,1,0,0,1,0,1,0,0,0,0,1,0,0,1,0,0,1,1,0,0,1,1,0,1,0},
            '{1,1,1,1,0,1,1,1,1,0,1,1,1,0,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,0,0,1,1,1,1,0,0,1,1,0,0,1,1,1,0,0,1,1,1,1,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,1,1,1,1,0,1,0,0,0,0,1,1,1,1,0,0,1,1,0,0,0,0,1,1,1,1,0,1,0,1,1,0,1,1,1,1,0,0,1,1,0,0,1,1,1,1,0},
            '{1,0,0,0,0,1,0,1,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,1,0,0,0,0,1,0,1,1,0,0,1,1,0,0,1,0,0,0,0,1,0,1,0,0,0,0,0,1,1,0,0,1,0,0,1,0,0,0,1,0,0,0,0,1,0,0,0,0,1,0,0,1,0,0,1,1,0,0,0,0,1,0,0,1,0,1,0,0,1,0,1,0,0,1,0,0,1,1,0,0,1,0,1,1,0},
            '{1,0,0,0,0,1,0,0,1,0,1,1,1,1,0,1,1,1,1,0,1,1,1,1,0,0,0,1,1,1,1,0,1,0,0,1,0,0,1,1,0,0,1,1,1,1,0,1,0,0,1,0,0,0,0,1,1,0,0,1,1,1,1,0,0,0,1,0,0,0,0,1,1,1,1,0,1,0,0,1,0,0,1,1,0,0,0,0,1,0,0,1,0,0,1,1,0,0,1,0,0,1,0,0,1,1,0,0,1,0,0,1,0}
        };
        
        high_score = '{
            '{5,0,0,5,0,0,5,5,0,0,0,5,5,0,0,5,0,0,5,0,0,0,5,5,5,5,0,0,5,5,5,0,0,5,5,0,0,5,5,5,5,0,5,5,5,5,0},
            '{5,0,0,5,0,0,5,5,0,0,5,0,0,0,0,5,0,0,5,0,0,0,5,0,0,0,0,5,0,0,0,0,5,0,0,5,0,5,0,0,5,0,5,0,0,0,0},
            '{5,5,5,5,0,0,5,5,0,0,5,0,5,5,0,5,5,5,5,0,0,0,5,5,5,5,0,5,0,0,0,0,5,0,0,5,0,5,5,5,5,0,5,5,5,0,0},
            '{5,0,0,5,0,0,5,5,0,0,5,0,0,5,0,5,0,0,5,0,0,0,0,0,0,5,0,5,0,0,0,0,5,0,0,5,0,5,0,5,0,0,5,0,0,0,0},
            '{5,0,0,5,0,0,5,5,0,0,0,5,5,0,0,5,0,0,5,0,0,0,5,5,5,5,0,0,5,5,5,0,0,5,5,0,0,5,0,0,5,0,5,5,5,5,0}
        };
        
        your_score = '{
            '{4,0,0,4,0,0,4,4,0,0,4,0,0,4,0,4,4,4,4,0,0,0,4,4,4,4,0,0,4,4,4,0,0,4,4,0,0,4,4,4,4,0,4,4,4,4,0},
            '{4,0,0,4,0,4,0,0,4,0,4,0,0,4,0,4,0,0,4,0,0,0,4,0,0,0,0,4,0,0,0,0,4,0,0,4,0,4,0,0,4,0,4,0,0,0,0},
            '{0,4,4,0,0,4,0,0,4,0,4,0,0,4,0,4,4,4,4,0,0,0,4,4,4,4,0,4,0,0,0,0,4,0,0,4,0,4,4,4,4,0,4,4,4,0,0},
            '{0,4,4,0,0,4,0,0,4,0,4,0,0,4,0,4,0,4,0,0,0,0,0,0,0,4,0,4,0,0,0,0,4,0,0,4,0,4,0,4,0,0,4,0,0,0,0},
            '{0,4,4,0,0,0,4,4,0,0,0,4,4,0,0,4,0,0,4,0,0,0,4,4,4,4,0,0,4,4,4,0,0,4,4,0,0,4,0,0,4,0,4,4,4,4,0}
        };
        
        score_letters = '{
            '{1,1,1,1,1,0,1,0,0,0,1,0,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1},
            '{0,0,0,0,1,0,0,1,0,0,1,0,1,0,0,0,1,0,0,0,0,0,1,0,1,0,0,0,0},
            '{1,1,1,1,1,0,1,1,1,1,1,0,1,0,0,0,1,0,0,0,0,0,1,0,1,1,1,1,1},
            '{0,0,0,0,1,0,1,0,0,0,1,0,1,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,1},
            '{1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1}
        };
		  
		level_letters = '{
			'{1,1,1,1,1,0,1,1,1,1,1,0,0,0,1,0,0,0,1,1,1,1,1,0,1,1,1,1,1},
            '{0,0,0,0,1,0,0,0,0,0,1,0,0,1,0,1,0,0,0,0,0,0,1,0,0,0,0,0,1},
            '{0,0,0,0,1,0,1,1,1,1,1,0,0,1,0,1,0,0,1,1,1,1,1,0,0,0,0,0,1},
            '{0,0,0,0,1,0,0,0,0,0,1,0,1,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,1},
            '{0,0,0,0,1,0,1,1,1,1,1,0,1,0,0,0,1,0,1,1,1,1,1,0,0,0,0,0,1}
        };
		  
		line_letters = '{
			'{1,1,1,1,1,0,1,0,0,0,1,0,0,0,1,0,0,0,1,1,1,1,1},
            '{0,0,0,0,1,0,1,1,0,0,1,0,0,0,1,0,0,0,0,0,0,0,1},
            '{1,1,1,1,1,0,1,0,1,0,1,0,0,0,1,0,0,0,0,0,0,0,1},
            '{0,0,0,0,1,0,1,0,0,1,1,0,0,0,1,0,0,0,0,0,0,0,1},
            '{1,1,1,1,1,0,1,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,1}
		  
		  };
            
        zero = '{
            '{9,9,9,9,9},
            '{9,0,0,0,9},
            '{9,0,0,0,9},
            '{9,0,0,0,9},
            '{9,9,9,9,9}
        };
            
            
        one = '{
            '{0,0,9,0,0},
            '{0,0,9,0,0},
            '{0,0,9,0,0},
            '{0,0,9,0,0},
            '{0,0,9,0,0}
        };	
            
        two = '{
            '{9,9,9,9,9},
            '{0,0,0,0,9},
            '{9,9,9,9,9},
            '{9,0,0,0,0},
            '{9,9,9,9,9}
        };

        three = '{
            '{9,9,9,9,9},
            '{9,0,0,0,0},
            '{9,9,9,9,9},
            '{9,0,0,0,0},
            '{9,9,9,9,9}
        };
            
            
            
        four = '{
            '{9,0,0,0,0},
            '{9,0,0,0,0},
            '{9,9,9,9,9},
            '{9,0,0,0,9},
            '{9,0,0,0,9}
        };
            
            
            
        five = '{
            '{9,9,9,9,9},
            '{9,0,0,0,0},
            '{9,9,9,9,9},
            '{0,0,0,0,9},
            '{9,9,9,9,9}
        };
            
            
            
            
        six = '{
            '{9,9,9,9,9},
            '{9,0,0,0,9},
            '{9,9,9,9,9},
            '{0,0,0,0,9},
            '{9,9,9,9,9}
        };
            
            
            
            
        seven = '{
            '{9,0,0,0,0},
            '{9,0,0,0,0},
            '{9,0,0,0,0},
            '{9,0,0,0,9},
            '{9,9,9,9,9}
        };

        eight = '{
            '{9,9,9,9,9},
            '{9,0,0,0,9},
            '{9,9,9,9,9},
            '{9,0,0,0,9},
            '{9,9,9,9,9}
        };	
            
        nine = '{
            '{9,9,9,9,9},
            '{9,0,0,0,0},
            '{9,9,9,9,9},
            '{9,0,0,0,9},
            '{9,9,9,9,9}
        };
        end
endmodule